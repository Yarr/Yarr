library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

package hw_type_pkg is
    constant c_HW_IDENT : std_logic_vector(7 downto 0) := x"04";
end hw_type_pkd;
